circuit
v1 0 n1 vac=5  vdc=0
L1 n1 n2 0.001
C1 n2 n3 0.0001
R1 n3 0 10
.end


















